----------------------------------------------------------------------------------
-- Company: TCD
-- Engineer: Brian Whelan
-- 
-- Create Date: 12.12.2020 20:42:53
-- Module Name: memory_32bit - Behavioral
-- Project Name: processor_project
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory_32bit is
 Port(
      address : in std_logic_vector(31 downto 0); 
      data_in : in std_logic_vector(31 downto 0);
      MW : in std_logic;
      Clk : in std_logic;
      data_out : out std_logic_vector(31 downto 0)
     );
end memory_32bit;

architecture Behavioral of memory_32bit is
    type mem_array is array(0 to 511) of std_logic_vector(31 downto 0);
begin
    mem_process : process(address, data_in, Clk)
        variable data_mem : mem_array := (
        --Data
        x"0000FFFF", x"FFFF0000", x"0000AAAA", x"AAAA0000",     --0 to 3    
        x"0000BBBB", x"BBBB0000", x"0000CCCC", x"CCCC0000",     --4 to 7    
        x"0000DDDD", x"DDDD0000", x"0000EEEE", x"EEEE0000",     --8 to 11   
        x"11111111", x"BBBBBBBB", x"00FFFF00", x"19334414",     --12 to 15
        
        x"00000000", x"00000000", x"00000000", x"00000000",     --16 to 19
        x"00000000", x"00000000", x"00000000", x"00000000",     --20 to 23
        x"00000000", x"00000000", x"00000000", x"00000000",     --24 to 27
        x"00000000", x"00000000", x"00000000", x"00000000",     --28 to 31
        x"00000000", x"00000000", x"00000000", x"00000000",     --32 to 35
        x"00000000", x"00000000", x"00000000", x"00000000",     --36 to 39
        x"00000000", x"00000000", x"00000000", x"00000000",     --40 to 43
        x"00000000", x"00000000", x"00000000", x"00000000",     --44 to 47
        x"00000000", x"00000000", x"00000000", x"00000000",     --48 to 51
        x"00000000", x"00000000", x"00000000", x"00000000",     --52 to 55
        x"00000000", x"00000000", x"00000000", x"00000000",     --56 to 59
        x"00000000", x"00000000", x"00000000", x"00000000",     --60 to 63  
        
        --Program/Instructions
        --                          Instruction             Pseudocode                      Opcode              DR    SA    SB     
        x"00008000",    --64        LD  R0, Memory[R0]      R0 = Memory[R0] = 0             00000000000000001   00000 00000 00000
        x"00008000",    --65        LD  R0, Memory[R0]      R0 = Memory[R0] = 0             00000000000000001   00000 00000 00000
        x"00008400",    --66        LD  R1, Memory[R0]      R1 = Memory[R0] = 0x0000FFFF    00000000000000001   00001 00000 00000
        x"00018000",    --67        INC R0, R0              R0 = R0 + 1 = 1                 00000000000000011   00000 00000 00000
        x"00008800",    --68        LD  R2, Memory[R0]      R2 = Memory[R0] = 0xFFFF0000    00000000000000001   00010 00000 00000
        x"00018000",    --69        INC R0, R0              R0 = R0 + 1 = 2                 00000000000000011   00000 00000 00000
        x"00008C00",    --70        LD  R3, Memory[R0]      R3 = Memory[R0] = 0x0000AAAA    00000000000000001   00011 00000 00000
        x"00018000",    --71        INC R0, R0              R0 = R0 + 1 = 3                 00000000000000011   00000 00000 00000
        x"00009000",    --72        LD  R4, Memory[R0]      R4 = Memory[R0] = 0xAAAA0000    00000000000000001   00100 00000 00000
        
        x"00001847",    --73        ADI R6, R2, #7          R6 = R2 + 7 = 0xFFFF0007        00000000000000000   00110 00010 00111
        x"0002A064",    --74        ADD R8, R3, R4          R8 = R3 + R4 = 0xAAAAAAAA       00000000000000101   01000 00011 00100
        x"00022900",    --75        NOT R10, R8             R10 = NOT R8 = 0x55555555       00000000000000100   01010 01000 00000
        x"00038802",    --76        SR  R2, R0, R2          R12 = (R2 >> R0) = 0x1FFFE000   00000000000000111   00010 00000 00010
        x"00060088",    --77  while CMP R4, R8              while(R4 != R8)                 00000000000001100   00000 00100 01000    
        x"00070004",    --78        BEQ stop                {                               00000000000001110   00000 00000 00100
        x"00029083",    --79        ADD R4, R4, R3              R4 = R4 + R3                00000000000000101   00100 00100 00011                                
        x"0006FC1B",    --80        B   while               }                               00000000000001101   11111 00000 11011
        x"00000000",    --81 
        x"0006FC1E",    --82  stop  B stop                                                  00000000000001101   11111 00000 11110  
        
        x"00000000",    --83     
        x"00000000",    --84 
        x"00000000",    --85 
        x"00000000",    --86 
        x"00000000",    --87     
        x"00000000",    --88 
        x"00000000",    --89 
        x"00000000",    --90 
        x"00000000",    --91    
        x"00000000",    --92 
        x"00000000",    --93 
        x"00000000",    --94 
        x"00000000",    --95   
        
        x"00000000", x"00000000", x"00000000", x"00000000",     --96 to 99
        x"00000000", x"00000000", x"00000000", x"00000000",     --100 to 103        
        x"00000000", x"00000000", x"00000000", x"00000000",     --104 to 107
        x"00000000", x"00000000", x"00000000", x"00000000",     --108 to 111
        x"00000000", x"00000000", x"00000000", x"00000000",     --112 to 115
        x"00000000", x"00000000", x"00000000", x"00000000",     --116 to 119
        x"00000000", x"00000000", x"00000000", x"00000000",     --120 to 123
        x"00000000", x"00000000", x"00000000", x"00000000",     --124 to 127
        x"00000000", x"00000000", x"00000000", x"00000000",     --128 to 131
        x"00000000", x"00000000", x"00000000", x"00000000",     --132 to 135
        x"00000000", x"00000000", x"00000000", x"00000000",     --136 to 139
        x"00000000", x"00000000", x"00000000", x"00000000",     --140 to 143
        x"00000000", x"00000000", x"00000000", x"00000000",     --144 to 147
        x"00000000", x"00000000", x"00000000", x"00000000",     --148 to 151
        x"00000000", x"00000000", x"00000000", x"00000000",     --152 to 155
        x"00000000", x"00000000", x"00000000", x"00000000",     --156 to 159
        x"00000000", x"00000000", x"00000000", x"00000000",     --160 to 163
        x"00000000", x"00000000", x"00000000", x"00000000",     --164 to 167
        x"00000000", x"00000000", x"00000000", x"00000000",     --168 to 171
        x"00000000", x"00000000", x"00000000", x"00000000",     --172 to 175
        x"00000000", x"00000000", x"00000000", x"00000000",     --176 to 179
        x"00000000", x"00000000", x"00000000", x"00000000",     --180 to 183
        x"00000000", x"00000000", x"00000000", x"00000000",     --184 to 187
        x"00000000", x"00000000", x"00000000", x"00000000",     --188 to 191
        x"00000000", x"00000000", x"00000000", x"00000000",     --192 to 195
        x"00000000", x"00000000", x"00000000", x"00000000",     --196 to 199
        x"00000000", x"00000000", x"00000000", x"00000000",     --200 to 203
        x"00000000", x"00000000", x"00000000", x"00000000",     --204 to 207
        x"00000000", x"00000000", x"00000000", x"00000000",     --208 to 211
        x"00000000", x"00000000", x"00000000", x"00000000",     --212 to 215
        x"00000000", x"00000000", x"00000000", x"00000000",     --216 to 219
        x"00000000", x"00000000", x"00000000", x"00000000",     --220 to 223
        x"00000000", x"00000000", x"00000000", x"00000000",     --224 to 227
        x"00000000", x"00000000", x"00000000", x"00000000",     --228 to 231
        x"00000000", x"00000000", x"00000000", x"00000000",     --232 to 235
        x"00000000", x"00000000", x"00000000", x"00000000",     --236 to 239
        x"00000000", x"00000000", x"00000000", x"00000000",     --240 to 243
        x"00000000", x"00000000", x"00000000", x"00000000",     --244 to 247
        x"00000000", x"00000000", x"00000000", x"00000000",     --248 to 251
        x"00000000", x"00000000", x"00000000", x"00000000",     --252 to 255
        x"00000000", x"00000000", x"00000000", x"00000000",     --256 to 259    
        x"00000000", x"00000000", x"00000000", x"00000000",     --260 to 263
        x"00000000", x"00000000", x"00000000", x"00000000",     --264 to 267
        x"00000000", x"00000000", x"00000000", x"00000000",     --268 to 271
        x"00000000", x"00000000", x"00000000", x"00000000",     --272 to 275
        x"00000000", x"00000000", x"00000000", x"00000000",     --276 to 279
        x"00000000", x"00000000", x"00000000", x"00000000",     --280 to 283
        x"00000000", x"00000000", x"00000000", x"00000000",     --284 to 287
        x"00000000", x"00000000", x"00000000", x"00000000",     --288 to 291
        x"00000000", x"00000000", x"00000000", x"00000000",     --292 to 295
        x"00000000", x"00000000", x"00000000", x"00000000",     --296 to 299
        x"00000000", x"00000000", x"00000000", x"00000000",     --300 to 303
        x"00000000", x"00000000", x"00000000", x"00000000",     --304 to 307
        x"00000000", x"00000000", x"00000000", x"00000000",     --308 to 311
        x"00000000", x"00000000", x"00000000", x"00000000",     --312 to 315
        x"00000000", x"00000000", x"00000000", x"00000000",     --316 to 319
        x"00000000", x"00000000", x"00000000", x"00000000",     --320 to 323
        x"00000000", x"00000000", x"00000000", x"00000000",     --324 to 327
        x"00000000", x"00000000", x"00000000", x"00000000",     --328 to 331
        x"00000000", x"00000000", x"00000000", x"00000000",     --332 to 335
        x"00000000", x"00000000", x"00000000", x"00000000",     --336 to 339
        x"00000000", x"00000000", x"00000000", x"00000000",     --340 to 343
        x"00000000", x"00000000", x"00000000", x"00000000",     --344 to 347
        x"00000000", x"00000000", x"00000000", x"00000000",     --348 to 351
        x"00000000", x"00000000", x"00000000", x"00000000",     --352 to 355
        x"00000000", x"00000000", x"00000000", x"00000000",     --356 to 359
        x"00000000", x"00000000", x"00000000", x"00000000",     --360 to 363
        x"00000000", x"00000000", x"00000000", x"00000000",     --364 to 367
        x"00000000", x"00000000", x"00000000", x"00000000",     --368 to 371
        x"00000000", x"00000000", x"00000000", x"00000000",     --372 to 375
        x"00000000", x"00000000", x"00000000", x"00000000",     --376 to 379
        x"00000000", x"00000000", x"00000000", x"00000000",     --380 to 383
        x"00000000", x"00000000", x"00000000", x"00000000",     --384 to 387
        x"00000000", x"00000000", x"00000000", x"00000000",     --388 to 391
        x"00000000", x"00000000", x"00000000", x"00000000",     --392 to 395
        x"00000000", x"00000000", x"00000000", x"00000000",     --396 to 399
        x"00000000", x"00000000", x"00000000", x"00000000",     --400 to 403
        x"00000000", x"00000000", x"00000000", x"00000000",     --404 to 407
        x"00000000", x"00000000", x"00000000", x"00000000",     --408 to 411
        x"00000000", x"00000000", x"00000000", x"00000000",     --412 to 415
        x"00000000", x"00000000", x"00000000", x"00000000",     --416 to 419
        x"00000000", x"00000000", x"00000000", x"00000000",     --420 to 423
        x"00000000", x"00000000", x"00000000", x"00000000",     --424 to 427
        x"00000000", x"00000000", x"00000000", x"00000000",     --428 to 431
        x"00000000", x"00000000", x"00000000", x"00000000",     --432 to 435
        x"00000000", x"00000000", x"00000000", x"00000000",     --436 to 439
        x"00000000", x"00000000", x"00000000", x"00000000",     --440 to 443
        x"00000000", x"00000000", x"00000000", x"00000000",     --444 to 447
        x"00000000", x"00000000", x"00000000", x"00000000",     --448 to 451
        x"00000000", x"00000000", x"00000000", x"00000000",     --452 to 455     
        x"00000000", x"00000000", x"00000000", x"00000000",     --456 to 459
        x"00000000", x"00000000", x"00000000", x"00000000",     --460 to 463
        x"00000000", x"00000000", x"00000000", x"00000000",     --464 to 467
        x"00000000", x"00000000", x"00000000", x"00000000",     --468 to 471
        x"00000000", x"00000000", x"00000000", x"00000000",     --472 to 475
        x"00000000", x"00000000", x"00000000", x"00000000",     --476 to 479
        x"00000000", x"00000000", x"00000000", x"00000000",     --480 to 483
        x"00000000", x"00000000", x"00000000", x"00000000",     --484 to 487
        x"00000000", x"00000000", x"00000000", x"00000000",     --488 to 491
        x"00000000", x"00000000", x"00000000", x"00000000",     --492 to 495
        x"00000000", x"00000000", x"00000000", x"00000000",     --496 to 499
        x"00000000", x"00000000", x"00000000", x"00000000",     --500 to 503
        x"00000000", x"00000000", x"00000000", x"00000000",     --504 to 507
        x"00000000", x"00000000", x"00000000", x"00000000");    --508 to 511
        variable addr : integer;
        begin
            addr := conv_integer(address(8 downto 0));
            if(MW = '1' AND Clk = '1') then
                data_mem(addr) := data_in;
            elsif(MW = '0' AND Clk = '1') then
                data_out <= data_mem(addr) after 5ns;
            end if;
    end process;
end Behavioral;
