----------------------------------------------------------------------------------
-- Company: TCD
-- Engineer: Brian Whelan
-- 
-- Create Date: 15.12.2020 10:05:54
-- Module Name: control_memory_32bit - Behavioral
-- Project Name: processor_project
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity control_memory_32bit is
 Port(
      in_CAR : in std_logic_vector(16 downto 0); 
      FL : out std_logic;                           -- 0
      RZ : out std_logic;                           -- 1
      RN : out std_logic;                           -- 2
      RC : out std_logic;                           -- 3
      RV : out std_logic;                           -- 4
      MW : out std_logic;                           -- 5
      MM : out std_logic;                           -- 6
      RW : out std_logic;                           -- 7
      MD : out std_logic;                           -- 8
      FS : out std_logic_vector(4 downto 0);        -- 9 to 13
      MB : out std_logic;                           -- 14
      TB : out std_logic;                           -- 15
      TA : out std_logic;                           -- 16
      TD : out std_logic;                           -- 17
      PL : out std_logic;                           -- 18
      PI : out std_logic;                           -- 19
      IL : out std_logic;                           -- 20
      MC : out std_logic;                           -- 21
      MS : out std_logic_vector(2 downto 0);        -- 22 to 24
      NA : out std_logic_vector(16 downto 0)        -- 25 to 41
     );
end control_memory_32bit;

architecture Behavioral of control_memory_32bit is
    type mem_array is array(0 to 255) of std_logic_vector(41 downto 0);
begin
    mem_process : process(in_CAR)
        variable control_mem : mem_array := (
--|41              25|24 22|21 |20 |19 |18 |17 |16 |15 |14 |13    9|8  |7  |6  |5  |4  |3  |2  |1  |0  |
--| Next Address(NA) | MS  |MC |IL |PI |PL |TD |TA |TB |MB |  FS   |MD |RW |MM |MW |RV |RC |RN |RZ |FL |
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"00010"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1", --00 (ADI)
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --01 (LD)
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0", --02 (ST)
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00001"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1", --03 (INC)
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01110"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1", --04 (NOT)
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00010"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1", --05 (ADD)
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --06 
  "00000000000001001"&"111"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"00000"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --07 (SR)
  "00000000000001001"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"10100"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --08 (SR shift)
  "00000000000001000"&"111"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"0"&"00110"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1", --09 (SR counter update)
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --0A (SR catch)
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --0B 
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"00101"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1", --0C (CMP)
  "00000000000010000"&"001"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --0D (B)
  "00000000000001101"&"100"&"0"&"0"&"0"&"0"&"1"&"1"&"1"&"0"&"00000"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --0E (BEQ)
  "00000000000010000"&"001"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --0F (BEQ catch)
  "00000000000010001"&"000"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0", --10 (Instruction Fetch)
  "00000000000000000"&"001"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --11 (Exit)
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --12
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --13
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --14
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --15
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --16 
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --17 
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --18
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --19
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --1A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --1B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --1C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --1D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --1E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --1F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --20 
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --21
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --22
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --23
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --24
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --25
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --26
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --27
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --28
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --29
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --2A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --2B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --2C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --2D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --2E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --2F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --30 
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --31
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --32
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --33
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --34
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --35
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --36
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --37
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --38
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --39
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --3A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --3B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --3C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --3D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --3E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --3F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --40 
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --41
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --42
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --43
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --44
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --45
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --46
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --47
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --48
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --49
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --4A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --4B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --4C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --4D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --4E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --4F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --50 
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --51
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --52
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --53
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --54
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --55
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --56
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --57
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --58
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --59
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --5A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --5B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --5C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --5D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --5E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --5F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --60 
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --61
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --62
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --63
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --64
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --65
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --66
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --67
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --68
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --69
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --6A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --6B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --6C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --6D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --6E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --6F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --70 
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --71
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --72
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --73
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --74
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --75
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --76
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --77
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --78
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --79
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --7A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --7B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --7C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --7D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --7E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --7F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --80
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --81
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --82
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --83
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --84
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --85
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --86
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --87
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --88
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --89
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --8A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --8B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --8C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --8D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --8E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --8F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --90
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --91
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --92
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --93
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --94
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --95
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --96
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --97
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --98
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --99
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --9A
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --9B
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --9C
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --9D
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --9E
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --9F
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A0
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A1
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A2
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A3
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A4
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A5
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A6
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A7
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A8
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --A9
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --AA
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --AB
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --AC
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --AD
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --AE
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --AF
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B0
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B1
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B2
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B3
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B4
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B5
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B6
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B7
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B8
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --B9
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --BA
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --BB
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --BC
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --BD
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --BE
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --BF
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C0
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C1
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C2
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C3
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C4
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C5
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C6
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C7
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C8
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --C9
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --CA
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --CB
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --CC
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --CD
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --CE
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --CF
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D0
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D1
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D2
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D3
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D4
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D5
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D6
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D7
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D8
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --D9
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --DA
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --DB
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --DC
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --DD
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --DE
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --DF
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E0
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E1
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E2
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E3
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E4
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E5
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E6
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E7
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E8
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --E9
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --EA
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --EB
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --EC
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --ED
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --EE
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --EF
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F0
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F1
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F2
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F3
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F4
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F5
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F6
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F7
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F8
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --F9
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --FA
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --FB
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --FC
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --FD
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0", --FE
  "00000000000000000"&"000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00000"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0");--FF
        variable addr : integer;
        variable control_out : std_logic_vector(41 downto 0);
        begin
            addr := conv_integer(in_CAR);
            control_out := control_mem(addr);
            FL <= control_out(0);
            RZ <= control_out(1);
            RN <= control_out(2);
            RC <= control_out(3);
            RV <= control_out(4);
            MW <= control_out(5);
            MM <= control_out(6);
            RW <= control_out(7);
            MD <= control_out(8);
            FS <= control_out(13 downto 9);
            MB <= control_out(14);
            TB <= control_out(15);
            TA <= control_out(16);
            TD <= control_out(17);
            PL <= control_out(18);
            PI <= control_out(19);
            IL <= control_out(20);
            MC <= control_out(21);
            MS <= control_out(24 downto 22);
            NA <= control_out(41 downto 25);
    end process;
end Behavioral;
